----------------------------------------------------------------------------------------------------
--    (c)2023 F. COLLIN
----------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.constants_pkg.all;

entity rom_start_screen is
    Port (
        clk : in std_logic;
        address : in std_logic_vector(12 downto 0); -- 6144 adresse (2^13 = 8192 < 6144)
        data : out std_logic_vector(RGB_LENGTH - 1 downto 0) -- color RVB 5-6-5
        );
end rom_start_screen;

architecture Behavioral of rom_start_screen is
    type rom_type is array (0 to 6143) of std_logic_vector(RGB_LENGTH - 1 downto 0);
    constant rom_data : rom_type := (
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0110011000101001",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "1111111100101100",
        "0110011000101001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0110011000101001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "1111111100101100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0110011000101001",
        "0110011000101001",
        "1111111100101100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0010001011101000",
        "0011110001001001",
        "0110011000101001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0110011000101001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0011110001001001",
        "0110011000101001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0110011000101001",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0011110001001001",
        "1111111100101100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0110011000101001",
        "0110011000101001",
        "1111111100101100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0110011000101001",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100111100111",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100111100111",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0010001011101000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0010001011101000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0110011000101001",
        "1111111100101100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0010001011101000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0010001011101000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0110011000101001",
        "0110011000101001",
        "0110011000101001",
        "0110011000101001",
        "1111111100101100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0110011000101001",
        "0110011000101001",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100111100111",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0110011000101001",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0011110001001001",
        "0011110001001001",
        "1111111100101100",
        "0110011000101001",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0110011000101001",
        "0110011000101001",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0110011000101001",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0110011000101001",
        "0110011000101001",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0110011000101001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0110011000101001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0110011000101001",
        "0001100010100100",
        "0010000101001000",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0110011000101001",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0110011000101001",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0110011000101001",
        "0110011000101001",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0001100111100111",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0010001011101000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0110011000101001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "1111111100101100",
        "0110011000101001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0010001011101000",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "1111111100101100",
        "0110011000101001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0010001011101000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0110011000101001",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0110011000101001",
        "0110011000101001",
        "0010001011101000",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0110011000101001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0110011000101001",
        "0110011000101001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100010100100",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0110011000101001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0110011000101001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0001100010100100",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0110011000101001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0110011000101001",
        "0110011000101001",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0001100111100111",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0110011000101001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0001100010100100",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0110011000101001",
        "0110011000101001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0110011000101001",
        "0011110001001001",
        "0011110001001001",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0001100010100100",
        "0001100111100111",
        "0011110001001001",
        "0001100111100111",
        "0001100111100111",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0010001011101000",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0011110001001001",
        "0110011000101001",
        "0001100010100100",
        "0110011000101001",
        "0011110001001001",
        "0011110001001001",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0011110001001001",
        "0011110001001001",
        "0001100111100111",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100111100111",
        "0011110001001001",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0110011000101001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100111100111",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0010001011101000",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0001100111100111",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0011110001001001",
        "0001100111100111",
        "0001100111100111",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0011110001001001",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0001100111100111",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0011110001001001",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0001100010100100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0001100010100100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010001011101000",
        "0010001011101000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0001100010100100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0010001011101000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0001100010100100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0001100010100100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0001100010100100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0001100010100100",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0011101000101100",
        "0011101000101100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0011101000101100",
        "0011101000101100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010001011101000",
        "0010001011101000",
        "0001100111100111",
        "0001100111100111",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0001100010100100",
        "0010000101001000",
        "0010000101001000",
        "0001100010100100",
        "0001100010100100",

    others => (others => '0')
    );
begin
                       
    process(clk, address)
    begin
        if rising_edge(clk) then
            data <= rom_data(to_integer(unsigned(address)));
        end if;
    end process;
                       
end Behavioral;
