library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity trans is
    port (
        nb_binaire : in std_logic_vector(7 downto 0); -- [0;255]
        s_cent, s_diz, s_unit : out std_logic_vector(6 downto 0)
    );
end trans;

architecture behav of trans is
begin
    process(nb_binaire)
    begin
        case (nb_binaire) is
            when "00000000" =>
                s_unit <= "0000001";
                s_diz <= "0000001";
                s_cent <= "0000001";
            
            when "00000001" =>
                s_unit <= "1001111";
                s_diz <= "0000001";
                s_cent <= "0000001";
            
            when "00000010" =>
                s_unit <= "0010010";
                s_diz <= "0000001";
                s_cent <= "0000001";
            
            when "00000011" =>
                s_unit <= "0000110";
                s_diz <= "0000001";
                s_cent <= "0000001";
            
            when "00000100" =>
                s_unit <= "1001100";
                s_diz <= "0000001";
                s_cent <= "0000001";
            
            when "00000101" =>
                s_unit <= "0100100";
                s_diz <= "0000001";
                s_cent <= "0000001";
            
            when "00000110" =>
                s_unit <= "0100000";
                s_diz <= "0000001";
                s_cent <= "0000001";
            
            when "00000111" =>
                s_unit <= "0001111";
                s_diz <= "0000001";
                s_cent <= "0000001";
            
            when "00001000" =>
                s_unit <= "0000000";
                s_diz <= "0000001";
                s_cent <= "0000001";
            
            when "00001001" =>
                s_unit <= "0000100";
                s_diz <= "0000001";
                s_cent <= "0000001";
            
            when "00001010" =>
                s_unit <= "0000001";
                s_diz <= "1001111";
                s_cent <= "0000001";
            
            when "00001011" =>
                s_unit <= "1001111";
                s_diz <= "1001111";
                s_cent <= "0000001";
            
            when "00001100" =>
                s_unit <= "0010010";
                s_diz <= "1001111";
                s_cent <= "0000001";
            
            when "00001101" =>
                s_unit <= "0000110";
                s_diz <= "1001111";
                s_cent <= "0000001";
            
            when "00001110" =>
                s_unit <= "1001100";
                s_diz <= "1001111";
                s_cent <= "0000001";
            
            when "00001111" =>
                s_unit <= "0100100";
                s_diz <= "1001111";
                s_cent <= "0000001";
            
            when "00010000" =>
                s_unit <= "0100000";
                s_diz <= "1001111";
                s_cent <= "0000001";
            
            when "00010001" =>
                s_unit <= "0001111";
                s_diz <= "1001111";
                s_cent <= "0000001";
            
            when "00010010" =>
                s_unit <= "0000000";
                s_diz <= "1001111";
                s_cent <= "0000001";
            
            when "00010011" =>
                s_unit <= "0000100";
                s_diz <= "1001111";
                s_cent <= "0000001";
            
            when "00010100" =>
                s_unit <= "0000001";
                s_diz <= "0010010";
                s_cent <= "0000001";
            
            when "00010101" =>
                s_unit <= "1001111";
                s_diz <= "0010010";
                s_cent <= "0000001";
            
            when "00010110" =>
                s_unit <= "0010010";
                s_diz <= "0010010";
                s_cent <= "0000001";
            
            when "00010111" =>
                s_unit <= "0000110";
                s_diz <= "0010010";
                s_cent <= "0000001";
            
            when "00011000" =>
                s_unit <= "1001100";
                s_diz <= "0010010";
                s_cent <= "0000001";
            
            when "00011001" =>
                s_unit <= "0100100";
                s_diz <= "0010010";
                s_cent <= "0000001";
            
            when "00011010" =>
                s_unit <= "0100000";
                s_diz <= "0010010";
                s_cent <= "0000001";
            
            when "00011011" =>
                s_unit <= "0001111";
                s_diz <= "0010010";
                s_cent <= "0000001";
            
            when "00011100" =>
                s_unit <= "0000000";
                s_diz <= "0010010";
                s_cent <= "0000001";
            
            when "00011101" =>
                s_unit <= "0000100";
                s_diz <= "0010010";
                s_cent <= "0000001";
            
            when "00011110" =>
                s_unit <= "0000001";
                s_diz <= "0000110";
                s_cent <= "0000001";
            
            when "00011111" =>
                s_unit <= "1001111";
                s_diz <= "0000110";
                s_cent <= "0000001";
            
            when "00100000" =>
                s_unit <= "0010010";
                s_diz <= "0000110";
                s_cent <= "0000001";
            
            when "00100001" =>
                s_unit <= "0000110";
                s_diz <= "0000110";
                s_cent <= "0000001";
            
            when "00100010" =>
                s_unit <= "1001100";
                s_diz <= "0000110";
                s_cent <= "0000001";
            
            when "00100011" =>
                s_unit <= "0100100";
                s_diz <= "0000110";
                s_cent <= "0000001";
            
            when "00100100" =>
                s_unit <= "0100000";
                s_diz <= "0000110";
                s_cent <= "0000001";
            
            when "00100101" =>
                s_unit <= "0001111";
                s_diz <= "0000110";
                s_cent <= "0000001";
            
            when "00100110" =>
                s_unit <= "0000000";
                s_diz <= "0000110";
                s_cent <= "0000001";
            
            when "00100111" =>
                s_unit <= "0000100";
                s_diz <= "0000110";
                s_cent <= "0000001";
            
            when "00101000" =>
                s_unit <= "0000001";
                s_diz <= "1001100";
                s_cent <= "0000001";
            
            when "00101001" =>
                s_unit <= "1001111";
                s_diz <= "1001100";
                s_cent <= "0000001";
            
            when "00101010" =>
                s_unit <= "0010010";
                s_diz <= "1001100";
                s_cent <= "0000001";
            
            when "00101011" =>
                s_unit <= "0000110";
                s_diz <= "1001100";
                s_cent <= "0000001";
            
            when "00101100" =>
                s_unit <= "1001100";
                s_diz <= "1001100";
                s_cent <= "0000001";
            
            when "00101101" =>
                s_unit <= "0100100";
                s_diz <= "1001100";
                s_cent <= "0000001";
            
            when "00101110" =>
                s_unit <= "0100000";
                s_diz <= "1001100";
                s_cent <= "0000001";
            
            when "00101111" =>
                s_unit <= "0001111";
                s_diz <= "1001100";
                s_cent <= "0000001";
            
            when "00110000" =>
                s_unit <= "0000000";
                s_diz <= "1001100";
                s_cent <= "0000001";
            
            when "00110001" =>
                s_unit <= "0000100";
                s_diz <= "1001100";
                s_cent <= "0000001";
            
            when "00110010" =>
                s_unit <= "0000001";
                s_diz <= "0100100";
                s_cent <= "0000001";
            
            when "00110011" =>
                s_unit <= "1001111";
                s_diz <= "0100100";
                s_cent <= "0000001";
            
            when "00110100" =>
                s_unit <= "0010010";
                s_diz <= "0100100";
                s_cent <= "0000001";
            
            when "00110101" =>
                s_unit <= "0000110";
                s_diz <= "0100100";
                s_cent <= "0000001";
            
            when "00110110" =>
                s_unit <= "1001100";
                s_diz <= "0100100";
                s_cent <= "0000001";
            
            when "00110111" =>
                s_unit <= "0100100";
                s_diz <= "0100100";
                s_cent <= "0000001";
            
            when "00111000" =>
                s_unit <= "0100000";
                s_diz <= "0100100";
                s_cent <= "0000001";
            
            when "00111001" =>
                s_unit <= "0001111";
                s_diz <= "0100100";
                s_cent <= "0000001";
            
            when "00111010" =>
                s_unit <= "0000000";
                s_diz <= "0100100";
                s_cent <= "0000001";
            
            when "00111011" =>
                s_unit <= "0000100";
                s_diz <= "0100100";
                s_cent <= "0000001";
            
            when "00111100" =>
                s_unit <= "0000001";
                s_diz <= "0100000";
                s_cent <= "0000001";
            
            when "00111101" =>
                s_unit <= "1001111";
                s_diz <= "0100000";
                s_cent <= "0000001";
            
            when "00111110" =>
                s_unit <= "0010010";
                s_diz <= "0100000";
                s_cent <= "0000001";
            
            when "00111111" =>
                s_unit <= "0000110";
                s_diz <= "0100000";
                s_cent <= "0000001";
            
            when "01000000" =>
                s_unit <= "1001100";
                s_diz <= "0100000";
                s_cent <= "0000001";
            
            when "01000001" =>
                s_unit <= "0100100";
                s_diz <= "0100000";
                s_cent <= "0000001";
            
            when "01000010" =>
                s_unit <= "0100000";
                s_diz <= "0100000";
                s_cent <= "0000001";
            
            when "01000011" =>
                s_unit <= "0001111";
                s_diz <= "0100000";
                s_cent <= "0000001";
            
            when "01000100" =>
                s_unit <= "0000000";
                s_diz <= "0100000";
                s_cent <= "0000001";
            
            when "01000101" =>
                s_unit <= "0000100";
                s_diz <= "0100000";
                s_cent <= "0000001";
            
            when "01000110" =>
                s_unit <= "0000001";
                s_diz <= "0001111";
                s_cent <= "0000001";
            
            when "01000111" =>
                s_unit <= "1001111";
                s_diz <= "0001111";
                s_cent <= "0000001";
            
            when "01001000" =>
                s_unit <= "0010010";
                s_diz <= "0001111";
                s_cent <= "0000001";
            
            when "01001001" =>
                s_unit <= "0000110";
                s_diz <= "0001111";
                s_cent <= "0000001";
            
            when "01001010" =>
                s_unit <= "1001100";
                s_diz <= "0001111";
                s_cent <= "0000001";
            
            when "01001011" =>
                s_unit <= "0100100";
                s_diz <= "0001111";
                s_cent <= "0000001";
            
            when "01001100" =>
                s_unit <= "0100000";
                s_diz <= "0001111";
                s_cent <= "0000001";
            
            when "01001101" =>
                s_unit <= "0001111";
                s_diz <= "0001111";
                s_cent <= "0000001";
            
            when "01001110" =>
                s_unit <= "0000000";
                s_diz <= "0001111";
                s_cent <= "0000001";
            
            when "01001111" =>
                s_unit <= "0000100";
                s_diz <= "0001111";
                s_cent <= "0000001";
            
            when "01010000" =>
                s_unit <= "0000001";
                s_diz <= "0000000";
                s_cent <= "0000001";
            
            when "01010001" =>
                s_unit <= "1001111";
                s_diz <= "0000000";
                s_cent <= "0000001";
            
            when "01010010" =>
                s_unit <= "0010010";
                s_diz <= "0000000";
                s_cent <= "0000001";
            
            when "01010011" =>
                s_unit <= "0000110";
                s_diz <= "0000000";
                s_cent <= "0000001";
            
            when "01010100" =>
                s_unit <= "1001100";
                s_diz <= "0000000";
                s_cent <= "0000001";
            
            when "01010101" =>
                s_unit <= "0100100";
                s_diz <= "0000000";
                s_cent <= "0000001";
            
            when "01010110" =>
                s_unit <= "0100000";
                s_diz <= "0000000";
                s_cent <= "0000001";
            
            when "01010111" =>
                s_unit <= "0001111";
                s_diz <= "0000000";
                s_cent <= "0000001";
            
            when "01011000" =>
                s_unit <= "0000000";
                s_diz <= "0000000";
                s_cent <= "0000001";
            
            when "01011001" =>
                s_unit <= "0000100";
                s_diz <= "0000000";
                s_cent <= "0000001";
            
            when "01011010" =>
                s_unit <= "0000001";
                s_diz <= "0000100";
                s_cent <= "0000001";
            
            when "01011011" =>
                s_unit <= "1001111";
                s_diz <= "0000100";
                s_cent <= "0000001";
            
            when "01011100" =>
                s_unit <= "0010010";
                s_diz <= "0000100";
                s_cent <= "0000001";
            
            when "01011101" =>
                s_unit <= "0000110";
                s_diz <= "0000100";
                s_cent <= "0000001";
            
            when "01011110" =>
                s_unit <= "1001100";
                s_diz <= "0000100";
                s_cent <= "0000001";
            
            when "01011111" =>
                s_unit <= "0100100";
                s_diz <= "0000100";
                s_cent <= "0000001";
            
            when "01100000" =>
                s_unit <= "0100000";
                s_diz <= "0000100";
                s_cent <= "0000001";
            
            when "01100001" =>
                s_unit <= "0001111";
                s_diz <= "0000100";
                s_cent <= "0000001";
            
            when "01100010" =>
                s_unit <= "0000000";
                s_diz <= "0000100";
                s_cent <= "0000001";
            
            when "01100011" =>
                s_unit <= "0000100";
                s_diz <= "0000100";
                s_cent <= "0000001";
            
            when "01100100" =>
                s_unit <= "0000001";
                s_diz <= "0000001";
                s_cent <= "1001111";
            
            when "01100101" =>
                s_unit <= "1001111";
                s_diz <= "0000001";
                s_cent <= "1001111";
            
            when "01100110" =>
                s_unit <= "0010010";
                s_diz <= "0000001";
                s_cent <= "1001111";
            
            when "01100111" =>
                s_unit <= "0000110";
                s_diz <= "0000001";
                s_cent <= "1001111";
            
            when "01101000" =>
                s_unit <= "1001100";
                s_diz <= "0000001";
                s_cent <= "1001111";
            
            when "01101001" =>
                s_unit <= "0100100";
                s_diz <= "0000001";
                s_cent <= "1001111";
            
            when "01101010" =>
                s_unit <= "0100000";
                s_diz <= "0000001";
                s_cent <= "1001111";
            
            when "01101011" =>
                s_unit <= "0001111";
                s_diz <= "0000001";
                s_cent <= "1001111";
            
            when "01101100" =>
                s_unit <= "0000000";
                s_diz <= "0000001";
                s_cent <= "1001111";
            
            when "01101101" =>
                s_unit <= "0000100";
                s_diz <= "0000001";
                s_cent <= "1001111";
            
            when "01101110" =>
                s_unit <= "0000001";
                s_diz <= "1001111";
                s_cent <= "1001111";
            
            when "01101111" =>
                s_unit <= "1001111";
                s_diz <= "1001111";
                s_cent <= "1001111";
            
            when "01110000" =>
                s_unit <= "0010010";
                s_diz <= "1001111";
                s_cent <= "1001111";
            
            when "01110001" =>
                s_unit <= "0000110";
                s_diz <= "1001111";
                s_cent <= "1001111";
            
            when "01110010" =>
                s_unit <= "1001100";
                s_diz <= "1001111";
                s_cent <= "1001111";
            
            when "01110011" =>
                s_unit <= "0100100";
                s_diz <= "1001111";
                s_cent <= "1001111";
            
            when "01110100" =>
                s_unit <= "0100000";
                s_diz <= "1001111";
                s_cent <= "1001111";
            
            when "01110101" =>
                s_unit <= "0001111";
                s_diz <= "1001111";
                s_cent <= "1001111";
            
            when "01110110" =>
                s_unit <= "0000000";
                s_diz <= "1001111";
                s_cent <= "1001111";
            
            when "01110111" =>
                s_unit <= "0000100";
                s_diz <= "1001111";
                s_cent <= "1001111";
            
            when "01111000" =>
                s_unit <= "0000001";
                s_diz <= "0010010";
                s_cent <= "1001111";
            
            when "01111001" =>
                s_unit <= "1001111";
                s_diz <= "0010010";
                s_cent <= "1001111";
            
            when "01111010" =>
                s_unit <= "0010010";
                s_diz <= "0010010";
                s_cent <= "1001111";
            
            when "01111011" =>
                s_unit <= "0000110";
                s_diz <= "0010010";
                s_cent <= "1001111";
            
            when "01111100" =>
                s_unit <= "1001100";
                s_diz <= "0010010";
                s_cent <= "1001111";
            
            when "01111101" =>
                s_unit <= "0100100";
                s_diz <= "0010010";
                s_cent <= "1001111";
            
            when "01111110" =>
                s_unit <= "0100000";
                s_diz <= "0010010";
                s_cent <= "1001111";
            
            when "01111111" =>
                s_unit <= "0001111";
                s_diz <= "0010010";
                s_cent <= "1001111";
            
            when "10000000" =>
                s_unit <= "0000000";
                s_diz <= "0010010";
                s_cent <= "1001111";
            
            when "10000001" =>
                s_unit <= "0000100";
                s_diz <= "0010010";
                s_cent <= "1001111";
            
            when "10000010" =>
                s_unit <= "0000001";
                s_diz <= "0000110";
                s_cent <= "1001111";
            
            when "10000011" =>
                s_unit <= "1001111";
                s_diz <= "0000110";
                s_cent <= "1001111";
            
            when "10000100" =>
                s_unit <= "0010010";
                s_diz <= "0000110";
                s_cent <= "1001111";
            
            when "10000101" =>
                s_unit <= "0000110";
                s_diz <= "0000110";
                s_cent <= "1001111";
            
            when "10000110" =>
                s_unit <= "1001100";
                s_diz <= "0000110";
                s_cent <= "1001111";
            
            when "10000111" =>
                s_unit <= "0100100";
                s_diz <= "0000110";
                s_cent <= "1001111";
            
            when "10001000" =>
                s_unit <= "0100000";
                s_diz <= "0000110";
                s_cent <= "1001111";
            
            when "10001001" =>
                s_unit <= "0001111";
                s_diz <= "0000110";
                s_cent <= "1001111";
            
            when "10001010" =>
                s_unit <= "0000000";
                s_diz <= "0000110";
                s_cent <= "1001111";
            
            when "10001011" =>
                s_unit <= "0000100";
                s_diz <= "0000110";
                s_cent <= "1001111";
            
            when "10001100" =>
                s_unit <= "0000001";
                s_diz <= "1001100";
                s_cent <= "1001111";
            
            when "10001101" =>
                s_unit <= "1001111";
                s_diz <= "1001100";
                s_cent <= "1001111";
            
            when "10001110" =>
                s_unit <= "0010010";
                s_diz <= "1001100";
                s_cent <= "1001111";
            
            when "10001111" =>
                s_unit <= "0000110";
                s_diz <= "1001100";
                s_cent <= "1001111";
            
            when "10010000" =>
                s_unit <= "1001100";
                s_diz <= "1001100";
                s_cent <= "1001111";
            
            when "10010001" =>
                s_unit <= "0100100";
                s_diz <= "1001100";
                s_cent <= "1001111";
            
            when "10010010" =>
                s_unit <= "0100000";
                s_diz <= "1001100";
                s_cent <= "1001111";
            
            when "10010011" =>
                s_unit <= "0001111";
                s_diz <= "1001100";
                s_cent <= "1001111";
            
            when "10010100" =>
                s_unit <= "0000000";
                s_diz <= "1001100";
                s_cent <= "1001111";
            
            when "10010101" =>
                s_unit <= "0000100";
                s_diz <= "1001100";
                s_cent <= "1001111";
            
            when "10010110" =>
                s_unit <= "0000001";
                s_diz <= "0100100";
                s_cent <= "1001111";
            
            when "10010111" =>
                s_unit <= "1001111";
                s_diz <= "0100100";
                s_cent <= "1001111";
            
            when "10011000" =>
                s_unit <= "0010010";
                s_diz <= "0100100";
                s_cent <= "1001111";
            
            when "10011001" =>
                s_unit <= "0000110";
                s_diz <= "0100100";
                s_cent <= "1001111";
            
            when "10011010" =>
                s_unit <= "1001100";
                s_diz <= "0100100";
                s_cent <= "1001111";
            
            when "10011011" =>
                s_unit <= "0100100";
                s_diz <= "0100100";
                s_cent <= "1001111";
            
            when "10011100" =>
                s_unit <= "0100000";
                s_diz <= "0100100";
                s_cent <= "1001111";
            
            when "10011101" =>
                s_unit <= "0001111";
                s_diz <= "0100100";
                s_cent <= "1001111";
            
            when "10011110" =>
                s_unit <= "0000000";
                s_diz <= "0100100";
                s_cent <= "1001111";
            
            when "10011111" =>
                s_unit <= "0000100";
                s_diz <= "0100100";
                s_cent <= "1001111";
            
            when "10100000" =>
                s_unit <= "0000001";
                s_diz <= "0100000";
                s_cent <= "1001111";
            
            when "10100001" =>
                s_unit <= "1001111";
                s_diz <= "0100000";
                s_cent <= "1001111";
            
            when "10100010" =>
                s_unit <= "0010010";
                s_diz <= "0100000";
                s_cent <= "1001111";
            
            when "10100011" =>
                s_unit <= "0000110";
                s_diz <= "0100000";
                s_cent <= "1001111";
            
            when "10100100" =>
                s_unit <= "1001100";
                s_diz <= "0100000";
                s_cent <= "1001111";
            
            when "10100101" =>
                s_unit <= "0100100";
                s_diz <= "0100000";
                s_cent <= "1001111";
            
            when "10100110" =>
                s_unit <= "0100000";
                s_diz <= "0100000";
                s_cent <= "1001111";
            
            when "10100111" =>
                s_unit <= "0001111";
                s_diz <= "0100000";
                s_cent <= "1001111";
            
            when "10101000" =>
                s_unit <= "0000000";
                s_diz <= "0100000";
                s_cent <= "1001111";
            
            when "10101001" =>
                s_unit <= "0000100";
                s_diz <= "0100000";
                s_cent <= "1001111";
            
            when "10101010" =>
                s_unit <= "0000001";
                s_diz <= "0001111";
                s_cent <= "1001111";
            
            when "10101011" =>
                s_unit <= "1001111";
                s_diz <= "0001111";
                s_cent <= "1001111";
            
            when "10101100" =>
                s_unit <= "0010010";
                s_diz <= "0001111";
                s_cent <= "1001111";
            
            when "10101101" =>
                s_unit <= "0000110";
                s_diz <= "0001111";
                s_cent <= "1001111";
            
            when "10101110" =>
                s_unit <= "1001100";
                s_diz <= "0001111";
                s_cent <= "1001111";
            
            when "10101111" =>
                s_unit <= "0100100";
                s_diz <= "0001111";
                s_cent <= "1001111";
            
            when "10110000" =>
                s_unit <= "0100000";
                s_diz <= "0001111";
                s_cent <= "1001111";
            
            when "10110001" =>
                s_unit <= "0001111";
                s_diz <= "0001111";
                s_cent <= "1001111";
            
            when "10110010" =>
                s_unit <= "0000000";
                s_diz <= "0001111";
                s_cent <= "1001111";
            
            when "10110011" =>
                s_unit <= "0000100";
                s_diz <= "0001111";
                s_cent <= "1001111";
            
            when "10110100" =>
                s_unit <= "0000001";
                s_diz <= "0000000";
                s_cent <= "1001111";
            
            when "10110101" =>
                s_unit <= "1001111";
                s_diz <= "0000000";
                s_cent <= "1001111";
            
            when "10110110" =>
                s_unit <= "0010010";
                s_diz <= "0000000";
                s_cent <= "1001111";
            
            when "10110111" =>
                s_unit <= "0000110";
                s_diz <= "0000000";
                s_cent <= "1001111";
            
            when "10111000" =>
                s_unit <= "1001100";
                s_diz <= "0000000";
                s_cent <= "1001111";
            
            when "10111001" =>
                s_unit <= "0100100";
                s_diz <= "0000000";
                s_cent <= "1001111";
            
            when "10111010" =>
                s_unit <= "0100000";
                s_diz <= "0000000";
                s_cent <= "1001111";
            
            when "10111011" =>
                s_unit <= "0001111";
                s_diz <= "0000000";
                s_cent <= "1001111";
            
            when "10111100" =>
                s_unit <= "0000000";
                s_diz <= "0000000";
                s_cent <= "1001111";
            
            when "10111101" =>
                s_unit <= "0000100";
                s_diz <= "0000000";
                s_cent <= "1001111";
            
            when "10111110" =>
                s_unit <= "0000001";
                s_diz <= "0000100";
                s_cent <= "1001111";
            
            when "10111111" =>
                s_unit <= "1001111";
                s_diz <= "0000100";
                s_cent <= "1001111";
            
            when "11000000" =>
                s_unit <= "0010010";
                s_diz <= "0000100";
                s_cent <= "1001111";
            
            when "11000001" =>
                s_unit <= "0000110";
                s_diz <= "0000100";
                s_cent <= "1001111";
            
            when "11000010" =>
                s_unit <= "1001100";
                s_diz <= "0000100";
                s_cent <= "1001111";
            
            when "11000011" =>
                s_unit <= "0100100";
                s_diz <= "0000100";
                s_cent <= "1001111";
            
            when "11000100" =>
                s_unit <= "0100000";
                s_diz <= "0000100";
                s_cent <= "1001111";
            
            when "11000101" =>
                s_unit <= "0001111";
                s_diz <= "0000100";
                s_cent <= "1001111";
            
            when "11000110" =>
                s_unit <= "0000000";
                s_diz <= "0000100";
                s_cent <= "1001111";
            
            when "11000111" =>
                s_unit <= "0000100";
                s_diz <= "0000100";
                s_cent <= "1001111";
            
            when "11001000" =>
                s_unit <= "0000001";
                s_diz <= "0000001";
                s_cent <= "0010010";
            
            when "11001001" =>
                s_unit <= "1001111";
                s_diz <= "0000001";
                s_cent <= "0010010";
            
            when "11001010" =>
                s_unit <= "0010010";
                s_diz <= "0000001";
                s_cent <= "0010010";
            
            when "11001011" =>
                s_unit <= "0000110";
                s_diz <= "0000001";
                s_cent <= "0010010";
            
            when "11001100" =>
                s_unit <= "1001100";
                s_diz <= "0000001";
                s_cent <= "0010010";
            
            when "11001101" =>
                s_unit <= "0100100";
                s_diz <= "0000001";
                s_cent <= "0010010";
            
            when "11001110" =>
                s_unit <= "0100000";
                s_diz <= "0000001";
                s_cent <= "0010010";
            
            when "11001111" =>
                s_unit <= "0001111";
                s_diz <= "0000001";
                s_cent <= "0010010";
            
            when "11010000" =>
                s_unit <= "0000000";
                s_diz <= "0000001";
                s_cent <= "0010010";
            
            when "11010001" =>
                s_unit <= "0000100";
                s_diz <= "0000001";
                s_cent <= "0010010";
            
            when "11010010" =>
                s_unit <= "0000001";
                s_diz <= "1001111";
                s_cent <= "0010010";
            
            when "11010011" =>
                s_unit <= "1001111";
                s_diz <= "1001111";
                s_cent <= "0010010";
            
            when "11010100" =>
                s_unit <= "0010010";
                s_diz <= "1001111";
                s_cent <= "0010010";
            
            when "11010101" =>
                s_unit <= "0000110";
                s_diz <= "1001111";
                s_cent <= "0010010";
            
            when "11010110" =>
                s_unit <= "1001100";
                s_diz <= "1001111";
                s_cent <= "0010010";
            
            when "11010111" =>
                s_unit <= "0100100";
                s_diz <= "1001111";
                s_cent <= "0010010";
            
            when "11011000" =>
                s_unit <= "0100000";
                s_diz <= "1001111";
                s_cent <= "0010010";
            
            when "11011001" =>
                s_unit <= "0001111";
                s_diz <= "1001111";
                s_cent <= "0010010";
            
            when "11011010" =>
                s_unit <= "0000000";
                s_diz <= "1001111";
                s_cent <= "0010010";
            
            when "11011011" =>
                s_unit <= "0000100";
                s_diz <= "1001111";
                s_cent <= "0010010";
            
            when "11011100" =>
                s_unit <= "0000001";
                s_diz <= "0010010";
                s_cent <= "0010010";
            
            when "11011101" =>
                s_unit <= "1001111";
                s_diz <= "0010010";
                s_cent <= "0010010";
            
            when "11011110" =>
                s_unit <= "0010010";
                s_diz <= "0010010";
                s_cent <= "0010010";
            
            when "11011111" =>
                s_unit <= "0000110";
                s_diz <= "0010010";
                s_cent <= "0010010";
            
            when "11100000" =>
                s_unit <= "1001100";
                s_diz <= "0010010";
                s_cent <= "0010010";
            
            when "11100001" =>
                s_unit <= "0100100";
                s_diz <= "0010010";
                s_cent <= "0010010";
            
            when "11100010" =>
                s_unit <= "0100000";
                s_diz <= "0010010";
                s_cent <= "0010010";
            
            when "11100011" =>
                s_unit <= "0001111";
                s_diz <= "0010010";
                s_cent <= "0010010";
            
            when "11100100" =>
                s_unit <= "0000000";
                s_diz <= "0010010";
                s_cent <= "0010010";
            
            when "11100101" =>
                s_unit <= "0000100";
                s_diz <= "0010010";
                s_cent <= "0010010";
            
            when "11100110" =>
                s_unit <= "0000001";
                s_diz <= "0000110";
                s_cent <= "0010010";
            
            when "11100111" =>
                s_unit <= "1001111";
                s_diz <= "0000110";
                s_cent <= "0010010";
            
            when "11101000" =>
                s_unit <= "0010010";
                s_diz <= "0000110";
                s_cent <= "0010010";
            
            when "11101001" =>
                s_unit <= "0000110";
                s_diz <= "0000110";
                s_cent <= "0010010";
            
            when "11101010" =>
                s_unit <= "1001100";
                s_diz <= "0000110";
                s_cent <= "0010010";
            
            when "11101011" =>
                s_unit <= "0100100";
                s_diz <= "0000110";
                s_cent <= "0010010";
            
            when "11101100" =>
                s_unit <= "0100000";
                s_diz <= "0000110";
                s_cent <= "0010010";
            
            when "11101101" =>
                s_unit <= "0001111";
                s_diz <= "0000110";
                s_cent <= "0010010";
            
            when "11101110" =>
                s_unit <= "0000000";
                s_diz <= "0000110";
                s_cent <= "0010010";
            
            when "11101111" =>
                s_unit <= "0000100";
                s_diz <= "0000110";
                s_cent <= "0010010";
            
            when "11110000" =>
                s_unit <= "0000001";
                s_diz <= "1001100";
                s_cent <= "0010010";
            
            when "11110001" =>
                s_unit <= "1001111";
                s_diz <= "1001100";
                s_cent <= "0010010";
            
            when "11110010" =>
                s_unit <= "0010010";
                s_diz <= "1001100";
                s_cent <= "0010010";
            
            when "11110011" =>
                s_unit <= "0000110";
                s_diz <= "1001100";
                s_cent <= "0010010";
            
            when "11110100" =>
                s_unit <= "1001100";
                s_diz <= "1001100";
                s_cent <= "0010010";
            
            when "11110101" =>
                s_unit <= "0100100";
                s_diz <= "1001100";
                s_cent <= "0010010";
            
            when "11110110" =>
                s_unit <= "0100000";
                s_diz <= "1001100";
                s_cent <= "0010010";
            
            when "11110111" =>
                s_unit <= "0001111";
                s_diz <= "1001100";
                s_cent <= "0010010";
            
            when "11111000" =>
                s_unit <= "0000000";
                s_diz <= "1001100";
                s_cent <= "0010010";
            
            when "11111001" =>
                s_unit <= "0000100";
                s_diz <= "1001100";
                s_cent <= "0010010";
            
            when "11111010" =>
                s_unit <= "0000001";
                s_diz <= "0100100";
                s_cent <= "0010010";
            
            when "11111011" =>
                s_unit <= "1001111";
                s_diz <= "0100100";
                s_cent <= "0010010";
            
            when "11111100" =>
                s_unit <= "0010010";
                s_diz <= "0100100";
                s_cent <= "0010010";
            
            when "11111101" =>
                s_unit <= "0000110";
                s_diz <= "0100100";
                s_cent <= "0010010";
            
            when "11111110" =>
                s_unit <= "1001100";
                s_diz <= "0100100";
                s_cent <= "0010010";
            
            when "11111111" =>
                s_unit <= "0100100";
                s_diz <= "0100100";
                s_cent <= "0010010";
            
            when others =>
                s_unit <= "0000100";
                s_diz <= "0000100";
                s_cent <= "0100100";
            end case;
    end process;  
end behav ;