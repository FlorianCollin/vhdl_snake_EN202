-- constants_pkg.vhdl
library ieee;
use ieee.std_logic_1164.all;

package constants_pkg is
  constant X_LENGTH : integer := 7;
  constant Y_LENGTH : integer := 6;
  constant RGB_LENGTH : integer := 16;
end package constants_pkg;

package body constants_pkg is
end package body constants_pkg;
